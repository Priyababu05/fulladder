module fulladder_gate_level
(input A,
 input B,
 input Cin,
 
 output S,
 output Cout );
        wire p,r,s;
               xor(p,A,B);
               xor(S,p,Cin);
               
               and(r,p,Cin);
               and(s,A,b);
               or(cout,r,s);
endmodule